BSV1    �&���  NST�  NFO    ��8d�  CPU 5  REG    ��{� 'RAM      3      � ��  ���       �       �                              �  H�    �    H��V    �V                                                H       �       �                                                                              �                           RYOUITI OOKUBO                                                                              �:ڑ����ɤ� �         � 2 PLAYERS�*�CONSTRUCTION�                                                                                          � H� @� H�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   FRM      CLK    ���	    APU 7  FRM    ��SQ0 5   REG       LEN     ENV      S00        @      SQ1 5   REG       LEN     ENV      S00        @      TRI &   REG        LEN     S00 	     !     NOI +   REG     LEN     ENV       S00    Y�@  DMC     REG    �     @    S00        DCB    S00                S00    O�  PPU W	  REG    ��    3PAL !    0<)	'  '8
;  OAM    � H� @� H�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   NMT                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ^k    00 HIk 20000                                                                               
               

                   
 
                                                                          

                    
  
                  
  
  
                                                                                                          1 PLAYER                                                        2 PLAYERS                                                       CONSTRUCTION                                                                                                                                                                                                                                                                                                                                         FRM    IMG �   MPR �   PRG    ACC    BNK              CHR *   ACC    BNK                     NMT    ACC    BNK              WRK    ACC    BNK       PRT    PD0     �PD1     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                